module char_decoder(
        output reg [255:0] OUT,
        input [2:0] IN
    );
    always @(*)
    begin
        case(IN[2:0])
                3'd1:  OUT = {{16{1'b0}}, {16{1'b0}}, {16{1'b0}}, 160'b0000000000100000_0000000000100000_0000000000100000_0000000000100000_0000000000100000_0000000000100000_0000000111100000_0000000000100000_0000000000100000_0000011111100000, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}}; // 'F'
                3'd2:  OUT = {{16{1'b0}}, {16{1'b0}}, {16{1'b0}}, 160'b0000011111100000_0000100000100000_0000100000100000_0000100000100000_0000100000100000_0000011111100000_0000001000100000_0000001000100000_0000001000100000_0000000111100000, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}}; // 'B'
                3'd3:  OUT = {{16{1'b0}}, {16{1'b0}}, {16{1'b0}}, 160'b0000001111000000_0000010000100000_0000010000000000_0000010000000000_0000010000000000_0000001111000000_0000000000100000_0000000000100000_0000010000100000_0000001111000000, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}}; // 'S'
                3'd4:  OUT = {{16{1'b0}}, {16{1'b0}}, {16{1'b0}}, 160'b0000011111100000_0000000000100000_0000000001000000_0000000010000000_0000000100000000_0000001000000000_0000010000000000_0000010000000000_0000010000100000_0000001111000000, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}}; // '2'
                3'd5:  OUT = {{16{1'b0}}, {16{1'b0}}, {16{1'b0}}, 160'b0000001111000000_0000010000100000_0000010000000000_0000010000000000_0000010000000000_0000001110000000_0000010000000000_0000010000000000_0000010000100000_0000001111000000, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}}; // '3'
                3'd6:  OUT = {{16{1'b0}}, {16{1'b0}}, {16{1'b0}}, 160'b0000000111000000_0000001000000000_0000010000000000_0000010000000000_0000011111000000_0000010000100000_0000010000100000_0000010000100000_0000010000100000_0000001111000000, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}}; // '9'
                3'd7:  OUT = {{16{1'b0}}, {16{1'b0}}, {16{1'b0}}, 160'b0000111100111000_0001000010010000_0001000010010000_0001000010010000_0001000010010000_0001000010010000_0001000010010000_0001000010010000_0001000010011000_0000111100010000, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}}; // '10'
                3'd8:  OUT = {{16{1'b0}}, {16{1'b0}}, {16{1'b0}}, 160'b0000000000100000_0000000000100000_0000000000100000_0000000000100000_0000000000100000_0000011111100000_0000010000100000_0000010000100000_0000010000100000_0000011111100000, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}}; // 'P'
                3'd9:  OUT = {{16{1'b0}}, {16{1'b0}}, {16{1'b0}}, 160'b0000000111000000_0000000010000000_0000000010000000_0000000010000000_0000000010000000_0000000010000000_0000000010000000_0000000010000000_0000000000110000_0000000010000000, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}}; // '1'
                3'd10: OUT = {{16{1'b0}}, {16{1'b0}}, {16{1'b0}}, 160'b0000111011100000_0001000100010000_0001000100010000_0001000100010000_0001000100010000_0001000000010000_0001000000010000_0001000000010000_0001000000010000_0001000000010000, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}}; // 'W'
                3'd11: OUT = {{16{1'b0}}, {16{1'b0}}, {16{1'b0}}, 160'b0000000111000000_0000000010000000_0000000010000000_0000000010000000_0000000010000000_0000000010000000_0000000010000000_0000000010000000_0000000010000000_0000000111000000, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}}; // 'I'
                3'd12: OUT = {{16{1'b0}}, {16{1'b0}}, {16{1'b0}}, 160'b0000010000100000_0000011000100000_0000011000100000_0000010100100000_0000010100100000_0000010010100000_0000010010100000_0000010001100000_0000010001100000_0000010000100000, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}}; // 'N'
                default: OUT = {256{1'b0}}; // empty
        endcase
    end
endmodule
